package Contexts;

import ModuleContext::*;
import ModuleCollect::*;

export ModuleContext::*;
export ModuleCollect::*;

endpackage
